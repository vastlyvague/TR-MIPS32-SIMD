`timescale 1ns / 1ps
/****************************** C E C S  4 4 0 ******************************
 * 
 * File Name:  BarrellShift_SIMD.v
 * Project:    Final_Project
 * Designer:   Thomas Nguyen and Reed Ellison
 * Email:      Tholinngu@gmail.com and notwreed@gmail.com
 * Rev. No.:   Version 1.0
 * Rev. Date:  04/20/2019
 *
 * Purpose: SIMD Barrel Shifter Module to shift vector content in registers.
 *
 * NoDes: 
 ****************************************************************************/
module BarrelShift_SIMD(simd_sel, D, type, shamt, Out);
   input [1:0] simd_sel;
   input       [4:0]   type;           // Function Select from MCU
   input       [4:0]   shamt;          // Shifting amount from IR[10:6]
   input      [31:0]   D;              // Data input for shifiDing
   output reg [31:0]   Out;            // Shifted Output
   
   always@(*)
      case(simd_sel)
      2'b01: //simd8
         case(type)
            5'h0E: // Shift Left Logical
               case(shamt)
                  5'd0:  Out = D;
                  5'd1:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[30:24], 1'b0}, {D[22:16], 1'b0},
                                {D[14:8],  1'b0}, {D[6:0],   1'b0}};
                  5'd2:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[29:24], 2'b0}, {D[21:16], 2'b0},
                                {D[13:8],  2'b0}, {D[5:0],   2'b0}};
                  5'd3:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[28:24], 3'b0}, {D[20:16], 3'b0},
                                {D[12:8],  3'b0}, {D[4:0],   3'b0}};
                  5'd4:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[27:24], 4'b0}, {D[19:16], 4'b0},
                                {D[11:8],  4'b0}, {D[3:0],   4'b0}};
                  5'd5:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[26:24], 5'b0}, {D[18:16], 5'b0},
                                {D[10:8],  5'b0}, {D[2:0],   5'b0}};
                  5'd6:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[25:24], 5'b0}, {D[17:16], 5'b0},
                                {D[9:8],   5'b0}, {D[1:0],   5'b0}};
                  5'd7:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[24], 6'b0}, {D[17], 6'b0},
                                {D[8],  6'b0}, {D[0],  6'b0}};
                  default: Out = 32'b0;
               endcase
            5'h0C: // Shift Right Logical
               case(shamt)
                  5'd0:  Out = D;
                  5'd1:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{1'b0, D[31:25]}, {1'b0, D[23:17]},
                                {1'b0, D[15:9]},  {1'b0, D[7:1]}};
                  5'd2:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{2'b0, D[31:26]}, {2'b0, D[23:18]},
                                {2'b0, D[15:10]}, {2'b0, D[7:2]}};
                  5'd3:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{3'b0, D[31:27]}, {3'b0, D[23:19]},
                                {3'b0, D[15:11]}, {3'b0, D[7:3]}};
                  5'd4:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{4'b0, D[31:28]}, {4'b0, D[23:20]},
                                {4'b0, D[15:12]}, {4'b0, D[7:4]}};
                  5'd5:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{5'b0, D[31:29]}, {5'b0, D[23:21]},
                                {5'b0, D[15:13]}, {5'b0, D[7:5]}};
                  5'd6:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{6'b0, D[31:30]}, {6'b0, D[23:22]},
                                {6'b0, D[15:14]}, {6'b0, D[7:6]}};
                  5'd7:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{7'b0, D[31]}, {7'b0, D[23]},
                                {7'b0, D[15]}, {7'b0, D[7]}};
                  default: Out = 32'b0;
               endcase
            5'h0D: // Shift Right Arithmetic
               case(shamt)
                  5'd0:  Out = D;
                  5'd1:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[31], D[31:25]}, {D[23], D[23:17]},
                                {D[15], D[15:9]},  {D[7], D[7:1]}};
                  5'd2:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{{2{D[31]}}, D[31:26]}, {{2{D[23]}}, D[23:18]},
                                {{2{D[15]}}, D[15:10]}, {{2{D[7]}}, D[7:2]}};
                  5'd3:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{{3{D[31]}}, D[31:27]}, {{3{D[23]}}, D[23:19]},
                                {{3{D[15]}}, D[15:11]}, {{3{D[7]}}, D[7:3]}};
                  5'd4:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{{4{D[31]}}, D[31:28]}, {{4{D[23]}}, D[23:20]},
                                {{4{D[15]}}, D[15:12]}, {{4{D[7]}}, D[7:4]}};
                  5'd5:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{{5{D[31]}}, D[31:29]}, {{5{D[23]}}, D[23:21]},
                                {{5{D[15]}}, D[15:13]}, {{5{D[7]}}, D[7:5]}};
                  5'd6:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{{6{D[31]}}, D[31:30]}, {{6{D[23]}}, D[23:22]},
                                {{6{D[15]}}, D[15:14]}, {{6{D[7]}}, D[7:6]}};
                  default:  Out = {{{7{D[31]}}, D[31]}, {{7{D[23]}}, D[23]},
                                  {{7{D[15]}}, D[15]},  {{7{D[7]}}, D[7]}};
               endcase
            5'h1A: // Rotate Left
               case(shamt)
                  5'd0:  Out = D;
                  5'd1:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[30:24], D[31]}, {D[22:16], D[23]},
                                {D[14:8],  D[15]}, {D[6:0],   D[7]}};
                  5'd2:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[29:24], D[31:30]}, {D[21:16], D[23:22]},
                                {D[13:8],  D[15:14]}, {D[5:0],   D[7:6]}};
                  5'd3:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[28:24], D[31:29]}, {D[20:16], D[23:21]},
                                {D[12:8],  D[15:13]}, {D[4:0],   D[7:5]}};
                  5'd4:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[27:24], D[31:28]}, {D[19:16], D[23:20]},
                                {D[11:8],  D[15:12]}, {D[3:0],   D[7:4]}};
                  5'd5:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[26:24], D[31:27]}, {D[18:16], D[23:19]},
                                {D[10:8],  D[15:11]}, {D[2:0],   D[7:3]}};
                  5'd6:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[25:24], D[31:26]}, {D[17:16], D[23:18]},
                                {D[9:8],   D[15:10]}, {D[1:0],   D[7:2]}};
                  5'd7:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[24], D[31:25]}, {D[16], D[23:17]},
                                {D[8],  D[15:9]},  {D[0],  D[7:1]}};
                  default: Out = D;
               endcase
            5'h1B: // Rotate Right
               case(shamt)
                  5'd0:  Out = D;
                  5'd1:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[24], D[31:25]}, {D[16], D[23:17]},
                                {D[8],  D[15:9]},  {D[0],  D[7:1]}};
                  5'd2:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[25:24], D[31:26]}, {D[17:16], D[23:18]},
                                {D[9:8],   D[15:10]}, {D[1:0],   D[7:2]}};
                  5'd3:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[26:24], D[31:27]}, {D[18:17], D[23:19]},
                                {D[10:8],  D[15:11]}, {D[2:0],   D[7:3]}};
                  5'd4:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[27:24], D[31:28]}, {D[19:17], D[23:20]},
                                {D[11:8],  D[15:12]}, {D[3:0],   D[7:4]}};
                  5'd5:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[28:24], D[31:29]}, {D[20:17], D[23:21]},
                                {D[12:8],  D[15:13]}, {D[4:0],   D[7:5]}};
                  5'd6:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[29:24], D[31:30]}, {D[21:17], D[23:22]},
                                {D[13:8],  D[15:14]}, {D[5:0],   D[7:6]}};
                  5'd7:  {Out[31:24], Out[23:16], Out[15:8], Out[7:0]}
                             = {{D[30:24], D[31]}, {D[22:17], D[23]},
                                {D[14:8],  D[15]}, {D[6:0],   D[7]}};
                  default: Out = D;
               endcase
         endcase
      2'b10: //simd16
         case(type)
            5'h0E: // Shift Left Logical
               case(shamt)     // 31:16 bits,            15:0 bits
                  5'd0:  Out = D;
                  5'd1:  {Out[31:16], Out[15:0]} =
                             {{D[30:16], 1'b0}, {D[14:0], 1'b0}};
                  5'd2:  {Out[31:16], Out[15:0]} =
                             {{D[29:16], 2'b0}, {D[13:0], 2'b0}};
                  5'd3:  {Out[31:16], Out[15:0]} =
                             {{D[28:16], 3'b0}, {D[12:0], 3'b0}};
                  5'd4:  {Out[31:16], Out[15:0]} =
                             {{D[27:16], 4'b0}, {D[11:0], 4'b0}};
                  5'd5:  {Out[31:16], Out[15:0]} =
                             {{D[26:16], 5'b0}, {D[10:0], 5'b0}};
                  5'd6:  {Out[31:16], Out[15:0]} =
                             {{D[25:16], 6'b0}, {D[9:0], 6'b0}};
                  5'd7:  {Out[31:16], Out[15:0]} =
                             {{D[24:16], 7'b0}, {D[8:0], 7'b0}};
                  5'd8:  {Out[31:16], Out[15:0]} =
                             {{D[23:16], 8'b0}, {D[7:0], 8'b0}};
                  5'd9:  {Out[31:16], Out[15:0]} =
                             {{D[22:16], 9'b0}, {D[6:0], 9'b0}};
                  5'd10:  {Out[31:16], Out[15:0]} =
                             {{D[21:16], 10'b0}, {D[5:0], 10'b0}};
                  5'd11:  {Out[31:16], Out[15:0]} =
                             {{D[20:16], 11'b0}, {D[4:0], 11'b0}};
                  5'd12:  {Out[31:16], Out[15:0]} =
                             {{D[19:16], 12'b0}, {D[3:0], 12'b0}};
                  5'd13:  {Out[31:16], Out[15:0]} =
                             {{D[18:16], 13'b0}, {D[2:0], 13'b0}};
                  5'd14:  {Out[31:16], Out[15:0]} =
                             {{D[17:16], 14'b0}, {D[1:0], 14'b0}};
                  5'd15:  {Out[31:16], Out[15:0]} =
                             {{D[16], 15'b0}, {D[0], 15'b0}};
                  default: Out = 32'b0;
               endcase
            5'h0C: // Shift Right Logical
               case(shamt)     // 31:16 bits,            15:0 bits
                  5'd0:  Out = D;
                  5'd1:  {Out[31:16],Out[15:0]} = 
                             {{1'b0, D[31:17]}, {1'b0, D[15:1]}};
                  5'd2:  {Out[31:16], Out[15:0]} =
                             {{2'b0, D[31:18]}, {2'b0, D[15:2]}};
                  5'd3:  {Out[31:16], Out[15:0]} =
                             {{3'b0, D[31:19]}, {3'b0, D[15:3]}};
                  5'd4:  {Out[31:16], Out[15:0]} =
                             {{4'b0, D[31:20]}, {4'b0, D[15:4]}};
                  5'd5:  {Out[31:16], Out[15:0]} =
                             {{5'b0, D[31:21]}, {5'b0, D[15:5]}};
                  5'd6:  {Out[31:16], Out[15:0]} =
                             {{6'b0, D[31:22]}, {6'b0, D[15:6]}};
                  5'd7:  {Out[31:16], Out[15:0]} =
                             {{7'b0, D[31:23]}, {7'b0, D[15:7]}};
                  5'd8:  {Out[31:16], Out[15:0]} =
                             {{8'b0, D[31:24]}, {8'b0, D[15:8]}};
                  5'd9:  {Out[31:16], Out[15:0]} =
                             {{9'b0, D[31:25]}, {9'b0, D[15:9]}};
                  5'd10:  {Out[31:16], Out[15:0]} =
                             {{10'b0, D[31:26]}, {10'b0, D[15:10]}};
                  5'd11:  {Out[31:16], Out[15:0]} =
                             {{11'b0, D[31:27]}, {11'b0, D[15:11]}};
                  5'd12:  {Out[31:16], Out[15:0]} =
                             {{12'b0, D[31:28]}, {12'b0, D[15:12]}};
                  5'd13:  {Out[31:16], Out[15:0]} =
                             {{13'b0, D[31:29]}, {13'b0, D[15:13]}};
                  5'd14:  {Out[31:16], Out[15:0]} =
                             {{14'b0, D[31:30]}, {14'b0, D[15:14]}};
                  5'd15:  {Out[31:16], Out[15:0]} =
                             {{15'b0, D[31]},    {15'b0, D[15]}};
                  default: Out = 32'b0;
               endcase
            5'h0D: // Shift Right Arithmetic
               case(shamt)     // 31:16 bits,            15:0 bits
                  5'd0:  Out = D;
                  5'd1:  {Out[31:16], Out[15:0]} =
                             {{{1{D[31]}}, D[31:17]}, {{1{D[15]}}, D[15:1]}};
                  5'd2:  {Out[31:16], Out[15:0]} =
                             {{{2{D[31]}}, D[31:18]}, {{2{D[15]}}, D[15:2]}};
                  5'd3:  {Out[31:16], Out[15:0]} =
                             {{{3{D[31]}}, D[31:19]}, {{3{D[15]}}, D[15:3]}};
                  5'd4:  {Out[31:16], Out[15:0]} =
                             {{{4{D[31]}}, D[31:20]}, {{4{D[15]}}, D[15:4]}};
                  5'd5:  {Out[31:16], Out[15:0]} =
                             {{{5{D[31]}}, D[31:21]}, {{5{D[15]}}, D[15:5]}};
                  5'd6:  {Out[31:16], Out[15:0]} =
                             {{{6{D[31]}}, D[31:22]}, {{6{D[15]}}, D[15:6]}};
                  5'd7:  {Out[31:16], Out[15:0]} =
                             {{{7{D[31]}}, D[31:23]}, {{7{D[15]}}, D[15:7]}};
                  5'd8:  {Out[31:16], Out[15:0]} =
                             {{{8{D[31]}}, D[31:24]}, {{8{D[15]}}, D[15:8]}};
                  5'd9:  {Out[31:16], Out[15:0]} =
                             {{{9{D[31]}}, D[31:25]}, {{9{D[15]}}, D[15:9]}};
                  5'd10:  {Out[31:16], Out[15:0]} =
                             {{{10{D[31]}}, D[31:26]}, {{10{D[15]}}, D[15:10]}};
                  5'd11:  {Out[31:16], Out[15:0]} =
                             {{{11{D[31]}}, D[31:27]}, {{11{D[15]}}, D[15:11]}};
                  5'd12:  {Out[31:16], Out[15:0]} =
                             {{{12{D[31]}}, D[31:28]}, {{12{D[15]}}, D[15:12]}};
                  5'd13:  {Out[31:16], Out[15:0]} =
                             {{{13{D[31]}}, D[31:29]}, {{13{D[15]}}, D[15:13]}};
                  5'd14:  {Out[31:16], Out[15:0]} =
                             {{{14{D[31]}}, D[31:30]}, {{14{D[15]}}, D[15:14]}};
                  5'd15:  {Out[31:16], Out[15:0]} =
                             {{{15{D[31]}}, D[31]},    {{15{D[15]}}, D[15]}};
                  default:  Out = {{16{D[31]}}, {16{D[15]}}};
               endcase
            5'h1A: // Rotate Left
               case(shamt)
                  5'd0:  Out = D;
                  5'd1:  {Out[31:16], Out[15:0]} =
                             {{D[30:16], D[31]},    {D[14:0], D[15]}};
                  5'd2:  {Out[31:16], Out[15:0]} =
                             {{D[29:16], D[31:30]}, {D[13:0], D[15:14]}};
                  5'd3:  {Out[31:16], Out[15:0]} =
                             {{D[28:16], D[31:29]}, {D[12:0], D[15:13]}};
                  5'd4:  {Out[31:16], Out[15:0]} =
                             {{D[27:16], D[31:28]}, {D[11:0], D[15:12]}};
                  5'd5:  {Out[31:16], Out[15:0]} =
                             {{D[26:16], D[31:27]}, {D[10:0], D[15:11]}};
                  5'd6:  {Out[31:16], Out[15:0]} =
                             {{D[25:16], D[31:26]}, {D[9:0],  D[15:10]}};
                  5'd7:  {Out[31:16], Out[15:0]} =
                             {{D[24:16], D[31:25]}, {D[8:0],  D[15:9]}};
                  5'd8:  {Out[31:16], Out[15:0]} =
                             {{D[23:16], D[31:24]}, {D[7:0],  D[15:8]}};
                  5'd9:  {Out[31:16], Out[15:0]} =
                             {{D[22:16], D[31:23]}, {D[6:0],  D[15:7]}};
                  5'd10:  {Out[31:16], Out[15:0]} =
                             {{D[21:16], D[31:22]}, {D[5:0], D[15:6]}};
                  5'd11:  {Out[31:16], Out[15:0]} =
                             {{D[20:16], D[31:21]}, {D[4:0], D[15:5]}};
                  5'd12:  {Out[31:16], Out[15:0]} =
                             {{D[19:16], D[31:20]}, {D[3:0], D[15:4]}};
                  5'd13:  {Out[31:16], Out[15:0]} =
                             {{D[18:16], D[31:19]}, {D[2:0], D[15:3]}};
                  5'd14:  {Out[31:16], Out[15:0]} =
                             {{D[17:16], D[31:18]}, {D[1:0], D[15:2]}};
                  5'd15:  {Out[31:16], Out[15:0]} =
                             {{D[16],    D[31:17]}, {D[0], D[15:1]}};
                  default: Out = D;
               endcase
            5'h1B: // Rotate Right
               case(shamt)
                  5'd0:  Out = D;
                  5'd1:  {Out[31:16], Out[15:0]} =
                             {{D[16], D[31:17]},    {D[0], D[15:1]}};
                  5'd2:  {Out[31:16], Out[15:0]} =
                             {{D[17:16], D[31:18]}, {D[1:0], D[15:2]}};
                  5'd3:  {Out[31:16], Out[15:0]} =
                             {{D[18:16], D[31:19]}, {D[2:0], D[15:3]}};
                  5'd4:  {Out[31:16], Out[15:0]} =
                             {{D[19:16], D[31:20]}, {D[3:0], D[15:4]}};
                  5'd5:  {Out[31:16], Out[15:0]} =
                             {{D[20:16], D[31:21]}, {D[4:0], D[15:5]}};
                  5'd6:  {Out[31:16], Out[15:0]} =
                             {{D[21:16], D[31:22]}, {D[5:0], D[15:6]}};
                  5'd7:  {Out[31:16], Out[15:0]} =
                             {{D[22:16], D[31:23]}, {D[6:0], D[15:7]}};
                  5'd8:  {Out[31:16], Out[15:0]} =
                             {{D[23:16], D[31:24]}, {D[7:0], D[15:8]}};
                  5'd9:  {Out[31:16], Out[15:0]} =
                             {{D[24:16], D[31:25]}, {D[8:0], D[15:9]}};
                  5'd10:  {Out[31:16], Out[15:0]} =
                             {{D[25:16], D[31:26]}, {D[9:0], D[15:10]}};
                  5'd11:  {Out[31:16], Out[15:0]} =
                             {{D[26:16], D[31:27]}, {D[10:0], D[15:11]}};
                  5'd12:  {Out[31:16], Out[15:0]} =
                             {{D[27:16], D[31:28]}, {D[11:0], D[15:12]}};
                  5'd13:  {Out[31:16], Out[15:0]} =
                             {{D[28:16], D[31:29]}, {D[12:0], D[15:13]}};
                  5'd14:  {Out[31:16], Out[15:0]} =
                             {{D[29:16], D[31:30]}, {D[13:0], D[15:14]}};
                  5'd15:  {Out[31:16], Out[15:0]} =
                             {{D[30:16], D[31]},    {D[14:0], D[15]}};
                  default: Out = D;
               endcase
         endcase
         default : Out = D;
      endcase
      
endmodule
