`timescale 1ns / 1ps
/****************************** C E C S  4 4 0 ******************************
 * 
 * File Name:  BarrellShifter.v
 * Project:    Final_Project
 * Designer:   Thomas Nguyen and Reed Ellison
 * Email:      Tholinngu@gmail.com and notwreed@gmail.com
 * Rev. No.:   Version 1.0
 * Rev. Date:  04/10/2019
 *
 * Purpose: Barrell Shifter Module Do Implement Dhe Shift Instructions
 * for the ALU
 *
 * NoDes: 
 ****************************************************************************/
module BarrellShifter(D, type, shamt, Out, C);
   
   input       [4:0]   type;           // Function Select from MCU
   input       [4:0]   shamt;          // Shifting amount from IR[10:6]
   input      [31:0]   D;              // Data input for shifiDing
   output reg          C;              // Carry flag
   output reg [31:0]   Out;            // Shifted Output
   
   always@(*)
      case(type)
         5'h0E: // Shift Left Logical
            case(shamt)
               5'd0:  {C,Out} = {1'b0, D};
               5'd1:  {C,Out} = {D[31], D[30:0],  1'b0};
               5'd2:  {C,Out} = {D[30], D[29:0],  2'b0};
               5'd3:  {C,Out} = {D[29], D[28:0],  3'b0};
               5'd4:  {C,Out} = {D[28], D[27:0],  4'b0};
               5'd5:  {C,Out} = {D[27], D[26:0],  5'b0};
               5'd6:  {C,Out} = {D[26], D[25:0],  6'b0};
               5'd7:  {C,Out} = {D[25], D[24:0],  7'b0};
               5'd8:  {C,Out} = {D[24], D[23:0],  8'b0};
               5'd9:  {C,Out} = {D[23], D[22:0],  9'b0};
               5'd10: {C,Out} = {D[22], D[21:0], 10'b0};
               5'd11: {C,Out} = {D[21], D[20:0], 11'b0};
               5'd12: {C,Out} = {D[20], D[19:0], 12'b0};
               5'd13: {C,Out} = {D[19], D[18:0], 13'b0};
               5'd14: {C,Out} = {D[18], D[17:0], 14'b0};
               5'd15: {C,Out} = {D[17], D[16:0], 15'b0};
               5'd16: {C,Out} = {D[16], D[15:0], 16'b0};
               5'd17: {C,Out} = {D[15], D[14:0], 17'b0};
               5'd18: {C,Out} = {D[14], D[13:0], 18'b0};
               5'd19: {C,Out} = {D[13], D[12:0], 19'b0};
               5'd20: {C,Out} = {D[12], D[11:0], 20'b0};
               5'd21: {C,Out} = {D[11], D[10:0], 21'b0};
               5'd22: {C,Out} = {D[10], D[ 9:0], 22'b0};
               5'd23: {C,Out} = {D[ 9], D[ 8:0], 23'b0};
               5'd24: {C,Out} = {D[ 8], D[ 7:0], 24'b0};
               5'd25: {C,Out} = {D[ 7], D[ 6:0], 25'b0};
               5'd26: {C,Out} = {D[ 6], D[ 5:0], 26'b0};
               5'd27: {C,Out} = {D[ 5], D[ 4:0], 27'b0};
               5'd28: {C,Out} = {D[ 4], D[ 3:0], 28'b0};
               5'd29: {C,Out} = {D[ 3], D[ 2:0], 29'b0};
               5'd30: {C,Out} = {D[ 2], D[ 1:0], 30'b0};
               5'd31: {C,Out} = {D[ 1], D[0],    31'b0};
            endcase
         5'h0C: // Shift Right Logical
            case(shamt)
               5'd0:  {C,Out} = {1'b0, D};
               5'd1:  {C,Out} = {D[ 0],  1'b0, D[31: 1]};
               5'd2:  {C,Out} = {D[ 1],  2'b0, D[31: 2]};
               5'd3:  {C,Out} = {D[ 2],  3'b0, D[31: 3]};
               5'd4:  {C,Out} = {D[ 3],  4'b0, D[31: 4]};
               5'd5:  {C,Out} = {D[ 4],  5'b0, D[31: 5]};
               5'd6:  {C,Out} = {D[ 5],  6'b0, D[31: 6]};
               5'd7:  {C,Out} = {D[ 6],  7'b0, D[31: 7]};
               5'd8:  {C,Out} = {D[ 7],  8'b0, D[31: 8]};
               5'd9:  {C,Out} = {D[ 8],  9'b0, D[31: 9]};
               5'd10: {C,Out} = {D[ 9], 10'b0, D[31:10]};
               5'd11: {C,Out} = {D[10], 11'b0, D[31:11]};
               5'd12: {C,Out} = {D[11], 12'b0, D[31:12]};
               5'd13: {C,Out} = {D[12], 13'b0, D[31:13]};
               5'd14: {C,Out} = {D[13], 14'b0, D[31:14]};
               5'd15: {C,Out} = {D[14], 15'b0, D[31:15]};
               5'd16: {C,Out} = {D[15], 16'b0, D[31:16]};
               5'd17: {C,Out} = {D[16], 17'b0, D[31:17]};
               5'd18: {C,Out} = {D[17], 18'b0, D[31:18]};
               5'd19: {C,Out} = {D[18], 19'b0, D[31:19]};
               5'd20: {C,Out} = {D[19], 20'b0, D[31:20]};
               5'd21: {C,Out} = {D[20], 21'b0, D[31:21]};
               5'd22: {C,Out} = {D[21], 22'b0, D[31:22]};
               5'd23: {C,Out} = {D[22], 23'b0, D[31:23]};
               5'd24: {C,Out} = {D[23], 24'b0, D[31:24]};
               5'd25: {C,Out} = {D[24], 25'b0, D[31:25]};
               5'd26: {C,Out} = {D[25], 26'b0, D[31:26]};
               5'd27: {C,Out} = {D[26], 27'b0, D[31:27]};
               5'd28: {C,Out} = {D[27], 28'b0, D[31:28]};
               5'd29: {C,Out} = {D[28], 29'b0, D[31:29]};
               5'd30: {C,Out} = {D[29], 30'b0, D[31:30]};
               5'd31: {C,Out} = {D[30], 31'b0, D[31]   };
            endcase
         5'h0D: // Shift Right Arithmetic
            case(shamt)
               5'd0:  {C,Out} = {1'b0, D};
               5'd1:  {C,Out} = {D[ 0], D[31], { 1{D[31]}}, D[30: 1]};
               5'd2:  {C,Out} = {D[ 1], D[31], { 2{D[31]}}, D[30: 2]};
               5'd3:  {C,Out} = {D[ 2], D[31], { 3{D[31]}}, D[30: 3]};
               5'd4:  {C,Out} = {D[ 3], D[31], { 4{D[31]}}, D[30: 4]};
               5'd5:  {C,Out} = {D[ 4], D[31], { 5{D[31]}}, D[30: 5]};
               5'd6:  {C,Out} = {D[ 5], D[31], { 6{D[31]}}, D[30: 6]};
               5'd7:  {C,Out} = {D[ 6], D[31], { 7{D[31]}}, D[30: 7]};
               5'd8:  {C,Out} = {D[ 7], D[31], { 8{D[31]}}, D[30: 8]};
               5'd9:  {C,Out} = {D[ 8], D[31], { 9{D[31]}}, D[30: 9]};
               5'd10: {C,Out} = {D[ 9], D[31], {10{D[31]}}, D[30:10]};
               5'd11: {C,Out} = {D[10], D[31], {11{D[31]}}, D[30:11]};
               5'd12: {C,Out} = {D[11], D[31], {12{D[31]}}, D[30:12]};
               5'd13: {C,Out} = {D[12], D[31], {13{D[31]}}, D[30:13]};
               5'd14: {C,Out} = {D[13], D[31], {14{D[31]}}, D[30:14]};
               5'd15: {C,Out} = {D[14], D[31], {15{D[31]}}, D[30:15]};
               5'd16: {C,Out} = {D[15], D[31], {16{D[31]}}, D[30:16]};
               5'd17: {C,Out} = {D[16], D[31], {17{D[31]}}, D[30:17]};
               5'd18: {C,Out} = {D[17], D[31], {18{D[31]}}, D[30:18]};
               5'd19: {C,Out} = {D[18], D[31], {19{D[31]}}, D[30:19]};
               5'd20: {C,Out} = {D[19], D[31], {20{D[31]}}, D[30:20]};
               5'd21: {C,Out} = {D[20], D[31], {21{D[31]}}, D[30:21]};
               5'd22: {C,Out} = {D[21], D[31], {22{D[31]}}, D[30:22]};
               5'd23: {C,Out} = {D[22], D[31], {23{D[31]}}, D[30:23]};
               5'd24: {C,Out} = {D[23], D[31], {24{D[31]}}, D[30:24]};
               5'd25: {C,Out} = {D[24], D[31], {25{D[31]}}, D[30:25]};
               5'd26: {C,Out} = {D[25], D[31], {26{D[31]}}, D[30:26]};
               5'd27: {C,Out} = {D[26], D[31], {27{D[31]}}, D[30:27]};
               5'd28: {C,Out} = {D[27], D[31], {28{D[31]}}, D[30:28]};
               5'd29: {C,Out} = {D[28], D[31], {29{D[31]}}, D[30:29]};
               5'd30: {C,Out} = {D[29], D[31], {30{D[31]}}, D[30]   };
               5'd31: {C,Out} = {D[30], D[31], {31{D[31]}}          };
            endcase
         5'h1A: // Rotate Left
            case(shamt)
               5'd0:  {C,Out} = D;
               5'd1:  {C,Out} = {D[30:0], D[31]};
               5'd2:  {C,Out} = {D[29:0], D[31:30]};
               5'd3:  {C,Out} = {D[28:0], D[31:29]};
               5'd4:  {C,Out} = {D[27:0], D[31:28]};
               5'd5:  {C,Out} = {D[26:0], D[31:27]};
               5'd6:  {C,Out} = {D[25:0], D[31:26]};
               5'd7:  {C,Out} = {D[24:0], D[31:25]};
               5'd8:  {C,Out} = {D[23:0], D[31:24]};
               5'd9:  {C,Out} = {D[22:0], D[31:23]};
               5'd10: {C,Out} = {D[21:0], D[31:22]};
               5'd11: {C,Out} = {D[20:0], D[31:21]};
               5'd12: {C,Out} = {D[19:0], D[31:20]};
               5'd13: {C,Out} = {D[18:0], D[31:19]};
               5'd14: {C,Out} = {D[17:0], D[31:18]};
               5'd15: {C,Out} = {D[16:0], D[31:17]};
               5'd16: {C,Out} = {D[15:0], D[31:16]};
               5'd17: {C,Out} = {D[14:0], D[31:15]};
               5'd18: {C,Out} = {D[13:0], D[31:14]};
               5'd19: {C,Out} = {D[12:0], D[31:13]};
               5'd20: {C,Out} = {D[11:0], D[31:12]};
               5'd21: {C,Out} = {D[10:0], D[31:11]};
               5'd22: {C,Out} = {D[9:0],  D[31:10]};
               5'd23: {C,Out} = {D[8:0],  D[31:9]};
               5'd24: {C,Out} = {D[7:0],  D[31:8]};
               5'd25: {C,Out} = {D[6:0],  D[31:7]};
               5'd26: {C,Out} = {D[5:0],  D[31:6]};
               5'd27: {C,Out} = {D[4:0],  D[31:5]};
               5'd28: {C,Out} = {D[3:0],  D[31:4]};
               5'd29: {C,Out} = {D[2:0],  D[31:3]};
               5'd30: {C,Out} = {D[1:0],  D[31:2]};
               5'd31: {C,Out} = {D[0],    D[31:1]};
            endcase
         5'h1B: // Rotate Right
            case(shamt)
               5'd0:  {C,Out} = D;
               5'd1:  {C,Out} = {D[0],    D[31:1]};
               5'd2:  {C,Out} = {D[1:0],  D[31:2]};
               5'd3:  {C,Out} = {D[2:0],  D[31:3]};
               5'd4:  {C,Out} = {D[3:0],  D[31:4]};
               5'd5:  {C,Out} = {D[4:0],  D[31:5]};
               5'd6:  {C,Out} = {D[5:0],  D[31:6]};
               5'd7:  {C,Out} = {D[6:0],  D[31:7]};
               5'd8:  {C,Out} = {D[7:0],  D[31:8]};
               5'd9:  {C,Out} = {D[8:0],  D[31:9]};
               5'd10: {C,Out} = {D[9:0],  D[31:10]};
               5'd11: {C,Out} = {D[10:0], D[31:11]};
               5'd12: {C,Out} = {D[11:0], D[31:12]};
               5'd13: {C,Out} = {D[12:0], D[31:13]};
               5'd14: {C,Out} = {D[13:0], D[31:14]};
               5'd15: {C,Out} = {D[14:0], D[31:15]};
               5'd16: {C,Out} = {D[15:0], D[31:16]};
               5'd17: {C,Out} = {D[16:0], D[31:17]};
               5'd18: {C,Out} = {D[17:0], D[31:18]};
               5'd19: {C,Out} = {D[18:0], D[31:19]};
               5'd20: {C,Out} = {D[19:0], D[31:20]};
               5'd21: {C,Out} = {D[20:0], D[31:21]};
               5'd22: {C,Out} = {D[21:0], D[31:22]};
               5'd23: {C,Out} = {D[22:0], D[31:23]};
               5'd24: {C,Out} = {D[23:0], D[31:24]};
               5'd25: {C,Out} = {D[24:0], D[31:25]};
               5'd26: {C,Out} = {D[25:0], D[31:26]};
               5'd27: {C,Out} = {D[26:0], D[31:27]};
               5'd28: {C,Out} = {D[27:0], D[31:28]};
               5'd29: {C,Out} = {D[28:0], D[31:29]};
               5'd30: {C,Out} = {D[29:0], D[31:30]};
               5'd31: {C,Out} = {D[30:0], D[31]};
            endcase
      endcase
      
endmodule
